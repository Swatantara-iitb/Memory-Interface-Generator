
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE ieee.numeric_std.ALL;


entity request_receive is
 port ( clk,rst: in std_logic;
        --ahir request interface
        ahir_request_req : in std_logic;
        ahir_request_ack : out std_logic;
        ahir_request_data: in std_logic_vector(63 downto 0);
       
      -- buffer interfaces 1 is for cmd_buf, 2 is for pend_buf
         wr_count1, wr_count2 : in integer range 0 to 9;
         wreq1, wreq2 : out std_logic;
         wack1, wack2 : in std_logic;
         wdata1, wdata2: out std_logic_vector(63 downto 0)
   
    );

end request_receive;  


architecture arch of request_receive is
 
--ahir data register 
component adr 
  port (clk, rst, adr_en : in std_logic;
        adr_in : in std_logic_vector(63 downto 0);
        adr_out: out std_logic_vector(63 downto 0)
       );

end component;

type state_type is (main, wait_on_1, wait_on_2, wait_on_count);
signal state: state_type;

signal flag : integer range 0 to 2;
-- adr interface
 
signal adr_en : std_logic;
signal adr_in, adr_out : std_logic_vector(63 downto 0);
   

-- command word parameters
signal cmd_check  : std_logic_vector(1 downto 0);
signal no_of_words  : integer range 0 to 8;
SIGNAL count_wr : INTEGER RANGE 0 TO 8 := 0;
signal rd_flag, wr_flag: integer range 0 to 1 := 0;


   begin 
      
   dut_adr : adr port map(clk, rst, adr_en, adr_in, adr_out);
    
      process(clk,state,rst)
        --variable words_count :integer range 0 to 8;
         begin
            if (rst = '1') then 
                state <= main;
            else if ( clk ='1' and clk 'event) then
                case state is
                      when main =>
                         flag <= 0; ahir_request_ack <= '0';
                        
                         -- request detected and count ok
                         if (ahir_request_req = '1' and wr_count1 <9 and wr_count2 < 9) then
                              wreq1 <= '1'; wreq2 <= '1'; flag <= 1 ;  
                             cmd_check <= ahir_request_data(63 downto 62);   
                             no_of_words <= to_integer(unsigned (ahir_request_data(55 downto 53))) ;
                             --words_count := no_of_words;
                              adr_en <= '1'; 
                              adr_in <= ahir_request_data;
                              -- read cmd
                              if (cmd_check = "00") then
                                rd_flag <= 1;
                              end if;
                             if (rd_flag = 1)  then
                                adr_en <= '1'; 
                                 if (wack1 = '1' and wack2 = '1' and ahir_request_req = '1' and wr_count1 <9 and wr_count2 <9   ) then

                                         wdata1 <= adr_out; wdata2 <= adr_out; adr_en <= '0';
                                         ahir_request_ack <= '1'; wreq1 <= '0'; wreq2 <= '0'; --rd_flag <= 0; 
                                 end if;
                                 
                             end if;
                             

                             -- write cmd
                             if (cmd_check = "01") then
                               wr_flag <= 1;
                             end if;
                             if (wr_flag = 1) then
                                      adr_en <= '1';
                                  if (wack1 = '1' and wack2 = '1' and ahir_request_req = '1'  ) then
                          
                                       if (count_wr <= (no_of_words+1) and wr_count1 <9 and wr_count2 <9 ) then
                                             adr_in <= ahir_request_data;
                                             wdata1 <= adr_out ; wdata2 <= adr_out;
                                             wreq1 <= '1'; wreq2 <= '1'; 
                                             count_wr <= count_wr + 1;
                                        else if (count_wr > no_of_words+1) then
                                             ahir_request_ack <= '1';
                                             wreq1 <= '0'; wreq2<= '0';
                                             adr_en <= '0';
                                                                                                                  
                                             end if;
                                       
                                        end if;
                                 
                                 end if;
                          
                            end if; 
                         end if;
                         -- count not ok
                         if ( ahir_request_req = '1' and (wr_count1 >9 or wr_count2 > 9) ) then
                              state <= wait_on_count;
                         end if;
                         
                         -- wait on 1
                         if (wack1 = '0' and wack2 = '1' and ahir_request_req = '1' and wr_count1 <9 and wr_count2 <9 ) then
                           wdata2 <= adr_out; wreq2 <= '0';
                           state <= wait_on_1;
                         end if;
                        
                         --wait on 2
                          if (wack1 = '1' and wack2 = '0' and ahir_request_req = '1' and wr_count1 <9 and wr_count2 <9 ) then
                             wdata1 <= adr_out; wreq1 <= '0';
                             state <= wait_on_2;
                          end if;                      




                      
                         
                      
                      
                    
            

                      when wait_on_1 =>
                         if (wack1 ='1' and ahir_request_req ='1' and wr_count1 <9  ) then
                             wdata1 <= adr_out;
                             ahir_request_ack <= '1';
                              wreq1 <= '0';
                              state <= main;

                        end if;
                         
                       when wait_on_2 =>
                         if (wack2 ='1' and ahir_request_req ='1' and wr_count2 <9 ) then
                             wdata2 <= adr_out;
                             ahir_request_ack <= '1';
                             wreq2 <= '0';
                              
                             state <= main;

                        end if;
                      
                    
                          
                        
                       when wait_on_count =>
                            if (wr_count1 <9 and wr_count2 <9 ) then
                               state <= main;
                                
                           end if;
                           if (flag = 0) then 
                               adr_en <= '1'; -- adr_en <= '1'; 
                               adr_in <= ahir_request_data;
                               ahir_request_ack <= '1';
                               flag <= 1;
                           end if;
                            if (flag = 1) then
                             adr_en <= '0'; 
                             end if;
                       end case;
                      end if;
                    end if;
                   end process;
end arch;    





                           

                             
        
